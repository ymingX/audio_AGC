// nios2.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module nios2 (
		input  wire        clk_clk,                                                //          clk.clk
		output wire [0:0]  flash_generic_tristate_controller_tcm_write_n_out,      //        flash.generic_tristate_controller_tcm_write_n_out
		output wire [0:0]  flash_generic_tristate_controller_tcm_chipselect_n_out, //             .generic_tristate_controller_tcm_chipselect_n_out
		output wire [0:0]  flash_generic_tristate_controller_tcm_read_n_out,       //             .generic_tristate_controller_tcm_read_n_out
		inout  wire [7:0]  flash_generic_tristate_controller_tcm_data_out,         //             .generic_tristate_controller_tcm_data_out
		output wire [21:0] flash_generic_tristate_controller_tcm_address_out,      //             .generic_tristate_controller_tcm_address_out
		input  wire [31:0] fmeasure_clk_export,                                    // fmeasure_clk.export
		input  wire [31:0] fmeasure_sqr_export,                                    // fmeasure_sqr.export
		input  wire [2:0]  keyirq_export,                                          //       keyirq.export
		input  wire [2:0]  keyvalue_export,                                        //     keyvalue.export
		output wire        lcd_lcd_cs_n,                                           //          lcd.lcd_cs_n
		output wire        lcd_lcd_wr_n,                                           //             .lcd_wr_n
		output wire        lcd_lcd_rd_n,                                           //             .lcd_rd_n
		output wire        lcd_lcd_rs,                                             //             .lcd_rs
		inout  wire [15:0] lcd_lcd_data,                                           //             .lcd_data
		input  wire        reset_reset_n,                                          //        reset.reset_n
		output wire [11:0] sdram_addr,                                             //        sdram.addr
		output wire [1:0]  sdram_ba,                                               //             .ba
		output wire        sdram_cas_n,                                            //             .cas_n
		output wire        sdram_cke,                                              //             .cke
		output wire        sdram_cs_n,                                             //             .cs_n
		inout  wire [15:0] sdram_dq,                                               //             .dq
		output wire [1:0]  sdram_dqm,                                              //             .dqm
		output wire        sdram_ras_n,                                            //             .ras_n
		output wire        sdram_we_n,                                             //             .we_n
		output wire        tas_scl_export,                                         //      tas_scl.export
		inout  wire        tas_sda_export,                                         //      tas_sda.export
		input  wire        touch_irq_export,                                       //    touch_irq.export
		output wire        touch_scl_export,                                       //    touch_scl.export
		inout  wire        touch_sda_export                                        //    touch_sda.export
	);

	wire         tristate_conduit_pin_sharer_tcm_request;                                              // tristate_conduit_pin_sharer:request -> tristate_conduit_bridge:request
	wire   [0:0] tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_read_n_out_out;       // tristate_conduit_pin_sharer:generic_tristate_controller_tcm_read_n_out -> tristate_conduit_bridge:tcs_generic_tristate_controller_tcm_read_n_out
	wire   [0:0] tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_write_n_out_out;      // tristate_conduit_pin_sharer:generic_tristate_controller_tcm_write_n_out -> tristate_conduit_bridge:tcs_generic_tristate_controller_tcm_write_n_out
	wire  [21:0] tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_address_out_out;      // tristate_conduit_pin_sharer:generic_tristate_controller_tcm_address_out -> tristate_conduit_bridge:tcs_generic_tristate_controller_tcm_address_out
	wire   [7:0] tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_data_out_out;         // tristate_conduit_pin_sharer:generic_tristate_controller_tcm_data_out -> tristate_conduit_bridge:tcs_generic_tristate_controller_tcm_data_out
	wire   [7:0] tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_data_out_in;          // tristate_conduit_bridge:tcs_generic_tristate_controller_tcm_data_in -> tristate_conduit_pin_sharer:generic_tristate_controller_tcm_data_in
	wire         tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_data_out_outen;       // tristate_conduit_pin_sharer:generic_tristate_controller_tcm_data_outen -> tristate_conduit_bridge:tcs_generic_tristate_controller_tcm_data_outen
	wire   [0:0] tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_chipselect_n_out_out; // tristate_conduit_pin_sharer:generic_tristate_controller_tcm_chipselect_n_out -> tristate_conduit_bridge:tcs_generic_tristate_controller_tcm_chipselect_n_out
	wire         tristate_conduit_pin_sharer_tcm_grant;                                                // tristate_conduit_bridge:grant -> tristate_conduit_pin_sharer:grant
	wire         generic_tristate_controller_tcm_data_outen;                                           // generic_tristate_controller:tcm_data_outen -> tristate_conduit_pin_sharer:tcs0_data_outen
	wire         generic_tristate_controller_tcm_request;                                              // generic_tristate_controller:tcm_request -> tristate_conduit_pin_sharer:tcs0_request
	wire         generic_tristate_controller_tcm_write_n_out;                                          // generic_tristate_controller:tcm_write_n_out -> tristate_conduit_pin_sharer:tcs0_write_n_out
	wire         generic_tristate_controller_tcm_read_n_out;                                           // generic_tristate_controller:tcm_read_n_out -> tristate_conduit_pin_sharer:tcs0_read_n_out
	wire         generic_tristate_controller_tcm_grant;                                                // tristate_conduit_pin_sharer:tcs0_grant -> generic_tristate_controller:tcm_grant
	wire         generic_tristate_controller_tcm_chipselect_n_out;                                     // generic_tristate_controller:tcm_chipselect_n_out -> tristate_conduit_pin_sharer:tcs0_chipselect_n_out
	wire  [21:0] generic_tristate_controller_tcm_address_out;                                          // generic_tristate_controller:tcm_address_out -> tristate_conduit_pin_sharer:tcs0_address_out
	wire   [7:0] generic_tristate_controller_tcm_data_out;                                             // generic_tristate_controller:tcm_data_out -> tristate_conduit_pin_sharer:tcs0_data_out
	wire   [7:0] generic_tristate_controller_tcm_data_in;                                              // tristate_conduit_pin_sharer:tcs0_data_in -> generic_tristate_controller:tcm_data_in
	wire  [31:0] cpu_data_master_readdata;                                                             // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                                          // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                                          // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [24:0] cpu_data_master_address;                                                              // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                                           // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                                                 // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                                                // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                                            // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                                                      // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                                                   // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [24:0] cpu_instruction_master_address;                                                       // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                                          // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                                                 // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                               // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                            // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                                   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                                  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_lcd_avalon_slave_chipselect;                                        // mm_interconnect_0:lcd_avalon_slave_chipselect -> lcd:cs_n
	wire  [31:0] mm_interconnect_0_lcd_avalon_slave_readdata;                                          // lcd:rddat -> mm_interconnect_0:lcd_avalon_slave_readdata
	wire   [0:0] mm_interconnect_0_lcd_avalon_slave_address;                                           // mm_interconnect_0:lcd_avalon_slave_address -> lcd:addr
	wire         mm_interconnect_0_lcd_avalon_slave_read;                                              // mm_interconnect_0:lcd_avalon_slave_read -> lcd:rd_n
	wire         mm_interconnect_0_lcd_avalon_slave_write;                                             // mm_interconnect_0:lcd_avalon_slave_write -> lcd:wr_n
	wire  [31:0] mm_interconnect_0_lcd_avalon_slave_writedata;                                         // mm_interconnect_0:lcd_avalon_slave_writedata -> lcd:wrdat
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                                       // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                                        // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;                                       // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;                                    // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;                                    // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;                                        // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                                           // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;                                     // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                                          // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;                                      // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_timer0_s1_chipselect;                                               // mm_interconnect_0:timer0_s1_chipselect -> timer0:chipselect
	wire  [15:0] mm_interconnect_0_timer0_s1_readdata;                                                 // timer0:readdata -> mm_interconnect_0:timer0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer0_s1_address;                                                  // mm_interconnect_0:timer0_s1_address -> timer0:address
	wire         mm_interconnect_0_timer0_s1_write;                                                    // mm_interconnect_0:timer0_s1_write -> timer0:write_n
	wire  [15:0] mm_interconnect_0_timer0_s1_writedata;                                                // mm_interconnect_0:timer0_s1_writedata -> timer0:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                                                // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                                  // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                               // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_s1_address;                                                   // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                                      // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                                // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                             // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                                     // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                                 // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_touch_irq_s1_chipselect;                                            // mm_interconnect_0:touch_irq_s1_chipselect -> touch_irq:chipselect
	wire  [31:0] mm_interconnect_0_touch_irq_s1_readdata;                                              // touch_irq:readdata -> mm_interconnect_0:touch_irq_s1_readdata
	wire   [1:0] mm_interconnect_0_touch_irq_s1_address;                                               // mm_interconnect_0:touch_irq_s1_address -> touch_irq:address
	wire         mm_interconnect_0_touch_irq_s1_write;                                                 // mm_interconnect_0:touch_irq_s1_write -> touch_irq:write_n
	wire  [31:0] mm_interconnect_0_touch_irq_s1_writedata;                                             // mm_interconnect_0:touch_irq_s1_writedata -> touch_irq:writedata
	wire         mm_interconnect_0_touch_sda_s1_chipselect;                                            // mm_interconnect_0:touch_sda_s1_chipselect -> touch_sda:chipselect
	wire  [31:0] mm_interconnect_0_touch_sda_s1_readdata;                                              // touch_sda:readdata -> mm_interconnect_0:touch_sda_s1_readdata
	wire   [1:0] mm_interconnect_0_touch_sda_s1_address;                                               // mm_interconnect_0:touch_sda_s1_address -> touch_sda:address
	wire         mm_interconnect_0_touch_sda_s1_write;                                                 // mm_interconnect_0:touch_sda_s1_write -> touch_sda:write_n
	wire  [31:0] mm_interconnect_0_touch_sda_s1_writedata;                                             // mm_interconnect_0:touch_sda_s1_writedata -> touch_sda:writedata
	wire         mm_interconnect_0_touch_scl_s1_chipselect;                                            // mm_interconnect_0:toucH_scl_s1_chipselect -> toucH_scl:chipselect
	wire  [31:0] mm_interconnect_0_touch_scl_s1_readdata;                                              // toucH_scl:readdata -> mm_interconnect_0:toucH_scl_s1_readdata
	wire   [1:0] mm_interconnect_0_touch_scl_s1_address;                                               // mm_interconnect_0:toucH_scl_s1_address -> toucH_scl:address
	wire         mm_interconnect_0_touch_scl_s1_write;                                                 // mm_interconnect_0:toucH_scl_s1_write -> toucH_scl:write_n
	wire  [31:0] mm_interconnect_0_touch_scl_s1_writedata;                                             // mm_interconnect_0:toucH_scl_s1_writedata -> toucH_scl:writedata
	wire         mm_interconnect_0_keyirq_s1_chipselect;                                               // mm_interconnect_0:keyirq_s1_chipselect -> keyirq:chipselect
	wire  [31:0] mm_interconnect_0_keyirq_s1_readdata;                                                 // keyirq:readdata -> mm_interconnect_0:keyirq_s1_readdata
	wire   [1:0] mm_interconnect_0_keyirq_s1_address;                                                  // mm_interconnect_0:keyirq_s1_address -> keyirq:address
	wire         mm_interconnect_0_keyirq_s1_write;                                                    // mm_interconnect_0:keyirq_s1_write -> keyirq:write_n
	wire  [31:0] mm_interconnect_0_keyirq_s1_writedata;                                                // mm_interconnect_0:keyirq_s1_writedata -> keyirq:writedata
	wire  [31:0] mm_interconnect_0_keyvalue_s1_readdata;                                               // keyvalue:readdata -> mm_interconnect_0:keyvalue_s1_readdata
	wire   [1:0] mm_interconnect_0_keyvalue_s1_address;                                                // mm_interconnect_0:keyvalue_s1_address -> keyvalue:address
	wire  [31:0] mm_interconnect_0_fmeasure_clk_s1_readdata;                                           // fmeasure_clk:readdata -> mm_interconnect_0:fmeasure_clk_s1_readdata
	wire   [1:0] mm_interconnect_0_fmeasure_clk_s1_address;                                            // mm_interconnect_0:fmeasure_clk_s1_address -> fmeasure_clk:address
	wire  [31:0] mm_interconnect_0_fmeasure_sqr_s1_readdata;                                           // fmeasure_sqr:readdata -> mm_interconnect_0:fmeasure_sqr_s1_readdata
	wire   [1:0] mm_interconnect_0_fmeasure_sqr_s1_address;                                            // mm_interconnect_0:fmeasure_sqr_s1_address -> fmeasure_sqr:address
	wire         mm_interconnect_0_tas_sda_s1_chipselect;                                              // mm_interconnect_0:TAS_sda_s1_chipselect -> TAS_sda:chipselect
	wire  [31:0] mm_interconnect_0_tas_sda_s1_readdata;                                                // TAS_sda:readdata -> mm_interconnect_0:TAS_sda_s1_readdata
	wire   [1:0] mm_interconnect_0_tas_sda_s1_address;                                                 // mm_interconnect_0:TAS_sda_s1_address -> TAS_sda:address
	wire         mm_interconnect_0_tas_sda_s1_write;                                                   // mm_interconnect_0:TAS_sda_s1_write -> TAS_sda:write_n
	wire  [31:0] mm_interconnect_0_tas_sda_s1_writedata;                                               // mm_interconnect_0:TAS_sda_s1_writedata -> TAS_sda:writedata
	wire         mm_interconnect_0_tas_scl_s1_chipselect;                                              // mm_interconnect_0:TAS_scl_s1_chipselect -> TAS_scl:chipselect
	wire  [31:0] mm_interconnect_0_tas_scl_s1_readdata;                                                // TAS_scl:readdata -> mm_interconnect_0:TAS_scl_s1_readdata
	wire   [1:0] mm_interconnect_0_tas_scl_s1_address;                                                 // mm_interconnect_0:TAS_scl_s1_address -> TAS_scl:address
	wire         mm_interconnect_0_tas_scl_s1_write;                                                   // mm_interconnect_0:TAS_scl_s1_write -> TAS_scl:write_n
	wire  [31:0] mm_interconnect_0_tas_scl_s1_writedata;                                               // mm_interconnect_0:TAS_scl_s1_writedata -> TAS_scl:writedata
	wire   [7:0] mm_interconnect_0_generic_tristate_controller_uas_readdata;                           // generic_tristate_controller:uas_readdata -> mm_interconnect_0:generic_tristate_controller_uas_readdata
	wire         mm_interconnect_0_generic_tristate_controller_uas_waitrequest;                        // generic_tristate_controller:uas_waitrequest -> mm_interconnect_0:generic_tristate_controller_uas_waitrequest
	wire         mm_interconnect_0_generic_tristate_controller_uas_debugaccess;                        // mm_interconnect_0:generic_tristate_controller_uas_debugaccess -> generic_tristate_controller:uas_debugaccess
	wire  [21:0] mm_interconnect_0_generic_tristate_controller_uas_address;                            // mm_interconnect_0:generic_tristate_controller_uas_address -> generic_tristate_controller:uas_address
	wire         mm_interconnect_0_generic_tristate_controller_uas_read;                               // mm_interconnect_0:generic_tristate_controller_uas_read -> generic_tristate_controller:uas_read
	wire   [0:0] mm_interconnect_0_generic_tristate_controller_uas_byteenable;                         // mm_interconnect_0:generic_tristate_controller_uas_byteenable -> generic_tristate_controller:uas_byteenable
	wire         mm_interconnect_0_generic_tristate_controller_uas_readdatavalid;                      // generic_tristate_controller:uas_readdatavalid -> mm_interconnect_0:generic_tristate_controller_uas_readdatavalid
	wire         mm_interconnect_0_generic_tristate_controller_uas_lock;                               // mm_interconnect_0:generic_tristate_controller_uas_lock -> generic_tristate_controller:uas_lock
	wire         mm_interconnect_0_generic_tristate_controller_uas_write;                              // mm_interconnect_0:generic_tristate_controller_uas_write -> generic_tristate_controller:uas_write
	wire   [7:0] mm_interconnect_0_generic_tristate_controller_uas_writedata;                          // mm_interconnect_0:generic_tristate_controller_uas_writedata -> generic_tristate_controller:uas_writedata
	wire   [0:0] mm_interconnect_0_generic_tristate_controller_uas_burstcount;                         // mm_interconnect_0:generic_tristate_controller_uas_burstcount -> generic_tristate_controller:uas_burstcount
	wire         irq_mapper_receiver0_irq;                                                             // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                             // timer0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                             // touch_irq:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                             // keyirq:irq -> irq_mapper:receiver3_irq
	wire  [31:0] cpu_irq_irq;                                                                          // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                                                       // rst_controller:reset_out -> [TAS_scl:reset_n, TAS_sda:reset_n, cpu:reset_n, fmeasure_clk:reset_n, fmeasure_sqr:reset_n, generic_tristate_controller:reset_reset, irq_mapper:reset, jtag_uart:rst_n, keyirq:reset_n, keyvalue:reset_n, lcd:rst_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram:reset_n, sysid:reset_n, timer0:reset_n, toucH_scl:reset_n, touch_irq:reset_n, touch_sda:reset_n, tristate_conduit_bridge:reset, tristate_conduit_pin_sharer:reset_reset]
	wire         rst_controller_reset_out_reset_req;                                                   // rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                                                        // cpu:debug_reset_request -> rst_controller:reset_in1

	nios2_TAS_scl tas_scl (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_tas_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tas_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tas_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tas_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tas_scl_s1_readdata),   //                    .readdata
		.out_port   (tas_scl_export)                           // external_connection.export
	);

	nios2_TAS_sda tas_sda (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_tas_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tas_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tas_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tas_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tas_sda_s1_readdata),   //                    .readdata
		.bidir_port (tas_sda_export)                           // external_connection.export
	);

	nios2_cpu cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	nios2_fmeasure_clk fmeasure_clk (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_fmeasure_clk_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_fmeasure_clk_s1_readdata), //                    .readdata
		.in_port  (fmeasure_clk_export)                         // external_connection.export
	);

	nios2_fmeasure_clk fmeasure_sqr (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_fmeasure_sqr_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_fmeasure_sqr_s1_readdata), //                    .readdata
		.in_port  (fmeasure_sqr_export)                         // external_connection.export
	);

	nios2_generic_tristate_controller #(
		.TCM_ADDRESS_W                  (22),
		.TCM_DATA_W                     (8),
		.TCM_BYTEENABLE_W               (1),
		.TCM_READ_WAIT                  (160),
		.TCM_WRITE_WAIT                 (160),
		.TCM_SETUP_WAIT                 (70),
		.TCM_DATA_HOLD                  (70),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (1),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) generic_tristate_controller (
		.clk_clk              (clk_clk),                                                         //   clk.clk
		.reset_reset          (rst_controller_reset_out_reset),                                  // reset.reset
		.uas_address          (mm_interconnect_0_generic_tristate_controller_uas_address),       //   uas.address
		.uas_burstcount       (mm_interconnect_0_generic_tristate_controller_uas_burstcount),    //      .burstcount
		.uas_read             (mm_interconnect_0_generic_tristate_controller_uas_read),          //      .read
		.uas_write            (mm_interconnect_0_generic_tristate_controller_uas_write),         //      .write
		.uas_waitrequest      (mm_interconnect_0_generic_tristate_controller_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (mm_interconnect_0_generic_tristate_controller_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable       (mm_interconnect_0_generic_tristate_controller_uas_byteenable),    //      .byteenable
		.uas_readdata         (mm_interconnect_0_generic_tristate_controller_uas_readdata),      //      .readdata
		.uas_writedata        (mm_interconnect_0_generic_tristate_controller_uas_writedata),     //      .writedata
		.uas_lock             (mm_interconnect_0_generic_tristate_controller_uas_lock),          //      .lock
		.uas_debugaccess      (mm_interconnect_0_generic_tristate_controller_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (generic_tristate_controller_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_read_n_out       (generic_tristate_controller_tcm_read_n_out),                      //      .read_n_out
		.tcm_chipselect_n_out (generic_tristate_controller_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_request          (generic_tristate_controller_tcm_request),                         //      .request
		.tcm_grant            (generic_tristate_controller_tcm_grant),                           //      .grant
		.tcm_address_out      (generic_tristate_controller_tcm_address_out),                     //      .address_out
		.tcm_data_out         (generic_tristate_controller_tcm_data_out),                        //      .data_out
		.tcm_data_outen       (generic_tristate_controller_tcm_data_outen),                      //      .data_outen
		.tcm_data_in          (generic_tristate_controller_tcm_data_in)                          //      .data_in
	);

	nios2_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	nios2_keyirq keyirq (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_keyirq_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keyirq_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keyirq_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keyirq_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keyirq_s1_readdata),   //                    .readdata
		.in_port    (keyirq_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                //                 irq.irq
	);

	nios2_keyvalue keyvalue (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_keyvalue_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_keyvalue_s1_readdata), //                    .readdata
		.in_port  (keyvalue_export)                         // external_connection.export
	);

	lcd lcd (
		.clk      (clk_clk),                                        //        clock.clk
		.wrdat    (mm_interconnect_0_lcd_avalon_slave_writedata),   // avalon_slave.writedata
		.rddat    (mm_interconnect_0_lcd_avalon_slave_readdata),    //             .readdata
		.cs_n     (~mm_interconnect_0_lcd_avalon_slave_chipselect), //             .chipselect_n
		.wr_n     (~mm_interconnect_0_lcd_avalon_slave_write),      //             .write_n
		.rd_n     (~mm_interconnect_0_lcd_avalon_slave_read),       //             .read_n
		.addr     (mm_interconnect_0_lcd_avalon_slave_address),     //             .address
		.lcd_cs_n (lcd_lcd_cs_n),                                   //  conduit_end.lcd_cs_n
		.lcd_wr_n (lcd_lcd_wr_n),                                   //             .lcd_wr_n
		.lcd_rd_n (lcd_lcd_rd_n),                                   //             .lcd_rd_n
		.lcd_rs   (lcd_lcd_rs),                                     //             .lcd_rs
		.lcd_data (lcd_lcd_data),                                   //             .lcd_data
		.rst_n    (~rst_controller_reset_out_reset)                 //        reset.reset_n
	);

	nios2_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	nios2_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	nios2_timer0 timer0 (
		.clk        (clk_clk),                                //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        // reset.reset_n
		.address    (mm_interconnect_0_timer0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                //   irq.irq
	);

	nios2_TAS_scl touch_scl (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_touch_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_touch_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_touch_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_touch_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_touch_scl_s1_readdata),   //                    .readdata
		.out_port   (touch_scl_export)                           // external_connection.export
	);

	nios2_touch_irq touch_irq (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_touch_irq_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_touch_irq_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_touch_irq_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_touch_irq_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_touch_irq_s1_readdata),   //                    .readdata
		.in_port    (touch_irq_export),                          // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                   //                 irq.irq
	);

	nios2_TAS_sda touch_sda (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_touch_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_touch_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_touch_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_touch_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_touch_sda_s1_readdata),   //                    .readdata
		.bidir_port (touch_sda_export)                           // external_connection.export
	);

	nios2_tristate_conduit_bridge tristate_conduit_bridge (
		.clk                                                  (clk_clk),                                                                              //   clk.clk
		.reset                                                (rst_controller_reset_out_reset),                                                       // reset.reset
		.request                                              (tristate_conduit_pin_sharer_tcm_request),                                              //   tcs.request
		.grant                                                (tristate_conduit_pin_sharer_tcm_grant),                                                //      .grant
		.tcs_generic_tristate_controller_tcm_write_n_out      (tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_write_n_out_out),      //      .generic_tristate_controller_tcm_write_n_out_out
		.tcs_generic_tristate_controller_tcm_chipselect_n_out (tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_chipselect_n_out_out), //      .generic_tristate_controller_tcm_chipselect_n_out_out
		.tcs_generic_tristate_controller_tcm_read_n_out       (tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_read_n_out_out),       //      .generic_tristate_controller_tcm_read_n_out_out
		.tcs_generic_tristate_controller_tcm_data_out         (tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_data_out_out),         //      .generic_tristate_controller_tcm_data_out_out
		.tcs_generic_tristate_controller_tcm_data_outen       (tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_data_out_outen),       //      .generic_tristate_controller_tcm_data_out_outen
		.tcs_generic_tristate_controller_tcm_data_in          (tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_data_out_in),          //      .generic_tristate_controller_tcm_data_out_in
		.tcs_generic_tristate_controller_tcm_address_out      (tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_address_out_out),      //      .generic_tristate_controller_tcm_address_out_out
		.generic_tristate_controller_tcm_write_n_out          (flash_generic_tristate_controller_tcm_write_n_out),                                    //   out.generic_tristate_controller_tcm_write_n_out
		.generic_tristate_controller_tcm_chipselect_n_out     (flash_generic_tristate_controller_tcm_chipselect_n_out),                               //      .generic_tristate_controller_tcm_chipselect_n_out
		.generic_tristate_controller_tcm_read_n_out           (flash_generic_tristate_controller_tcm_read_n_out),                                     //      .generic_tristate_controller_tcm_read_n_out
		.generic_tristate_controller_tcm_data_out             (flash_generic_tristate_controller_tcm_data_out),                                       //      .generic_tristate_controller_tcm_data_out
		.generic_tristate_controller_tcm_address_out          (flash_generic_tristate_controller_tcm_address_out)                                     //      .generic_tristate_controller_tcm_address_out
	);

	nios2_tristate_conduit_pin_sharer tristate_conduit_pin_sharer (
		.clk_clk                                          (clk_clk),                                                                              //   clk.clk
		.reset_reset                                      (rst_controller_reset_out_reset),                                                       // reset.reset
		.request                                          (tristate_conduit_pin_sharer_tcm_request),                                              //   tcm.request
		.grant                                            (tristate_conduit_pin_sharer_tcm_grant),                                                //      .grant
		.generic_tristate_controller_tcm_address_out      (tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_address_out_out),      //      .generic_tristate_controller_tcm_address_out_out
		.generic_tristate_controller_tcm_read_n_out       (tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_read_n_out_out),       //      .generic_tristate_controller_tcm_read_n_out_out
		.generic_tristate_controller_tcm_write_n_out      (tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_write_n_out_out),      //      .generic_tristate_controller_tcm_write_n_out_out
		.generic_tristate_controller_tcm_data_out         (tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_data_out_out),         //      .generic_tristate_controller_tcm_data_out_out
		.generic_tristate_controller_tcm_data_in          (tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_data_out_in),          //      .generic_tristate_controller_tcm_data_out_in
		.generic_tristate_controller_tcm_data_outen       (tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_data_out_outen),       //      .generic_tristate_controller_tcm_data_out_outen
		.generic_tristate_controller_tcm_chipselect_n_out (tristate_conduit_pin_sharer_tcm_generic_tristate_controller_tcm_chipselect_n_out_out), //      .generic_tristate_controller_tcm_chipselect_n_out_out
		.tcs0_request                                     (generic_tristate_controller_tcm_request),                                              //  tcs0.request
		.tcs0_grant                                       (generic_tristate_controller_tcm_grant),                                                //      .grant
		.tcs0_address_out                                 (generic_tristate_controller_tcm_address_out),                                          //      .address_out
		.tcs0_read_n_out                                  (generic_tristate_controller_tcm_read_n_out),                                           //      .read_n_out
		.tcs0_write_n_out                                 (generic_tristate_controller_tcm_write_n_out),                                          //      .write_n_out
		.tcs0_data_out                                    (generic_tristate_controller_tcm_data_out),                                             //      .data_out
		.tcs0_data_in                                     (generic_tristate_controller_tcm_data_in),                                              //      .data_in
		.tcs0_data_outen                                  (generic_tristate_controller_tcm_data_outen),                                           //      .data_outen
		.tcs0_chipselect_n_out                            (generic_tristate_controller_tcm_chipselect_n_out)                                      //      .chipselect_n_out
	);

	nios2_mm_interconnect_0 mm_interconnect_0 (
		.clk_100M_clk_clk                              (clk_clk),                                                         //                    clk_100M_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                                  // cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                       (cpu_data_master_address),                                         //                 cpu_data_master.address
		.cpu_data_master_waitrequest                   (cpu_data_master_waitrequest),                                     //                                .waitrequest
		.cpu_data_master_byteenable                    (cpu_data_master_byteenable),                                      //                                .byteenable
		.cpu_data_master_read                          (cpu_data_master_read),                                            //                                .read
		.cpu_data_master_readdata                      (cpu_data_master_readdata),                                        //                                .readdata
		.cpu_data_master_write                         (cpu_data_master_write),                                           //                                .write
		.cpu_data_master_writedata                     (cpu_data_master_writedata),                                       //                                .writedata
		.cpu_data_master_debugaccess                   (cpu_data_master_debugaccess),                                     //                                .debugaccess
		.cpu_instruction_master_address                (cpu_instruction_master_address),                                  //          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest            (cpu_instruction_master_waitrequest),                              //                                .waitrequest
		.cpu_instruction_master_read                   (cpu_instruction_master_read),                                     //                                .read
		.cpu_instruction_master_readdata               (cpu_instruction_master_readdata),                                 //                                .readdata
		.cpu_instruction_master_readdatavalid          (cpu_instruction_master_readdatavalid),                            //                                .readdatavalid
		.cpu_debug_mem_slave_address                   (mm_interconnect_0_cpu_debug_mem_slave_address),                   //             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                     (mm_interconnect_0_cpu_debug_mem_slave_write),                     //                                .write
		.cpu_debug_mem_slave_read                      (mm_interconnect_0_cpu_debug_mem_slave_read),                      //                                .read
		.cpu_debug_mem_slave_readdata                  (mm_interconnect_0_cpu_debug_mem_slave_readdata),                  //                                .readdata
		.cpu_debug_mem_slave_writedata                 (mm_interconnect_0_cpu_debug_mem_slave_writedata),                 //                                .writedata
		.cpu_debug_mem_slave_byteenable                (mm_interconnect_0_cpu_debug_mem_slave_byteenable),                //                                .byteenable
		.cpu_debug_mem_slave_waitrequest               (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),               //                                .waitrequest
		.cpu_debug_mem_slave_debugaccess               (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),               //                                .debugaccess
		.fmeasure_clk_s1_address                       (mm_interconnect_0_fmeasure_clk_s1_address),                       //                 fmeasure_clk_s1.address
		.fmeasure_clk_s1_readdata                      (mm_interconnect_0_fmeasure_clk_s1_readdata),                      //                                .readdata
		.fmeasure_sqr_s1_address                       (mm_interconnect_0_fmeasure_sqr_s1_address),                       //                 fmeasure_sqr_s1.address
		.fmeasure_sqr_s1_readdata                      (mm_interconnect_0_fmeasure_sqr_s1_readdata),                      //                                .readdata
		.generic_tristate_controller_uas_address       (mm_interconnect_0_generic_tristate_controller_uas_address),       // generic_tristate_controller_uas.address
		.generic_tristate_controller_uas_write         (mm_interconnect_0_generic_tristate_controller_uas_write),         //                                .write
		.generic_tristate_controller_uas_read          (mm_interconnect_0_generic_tristate_controller_uas_read),          //                                .read
		.generic_tristate_controller_uas_readdata      (mm_interconnect_0_generic_tristate_controller_uas_readdata),      //                                .readdata
		.generic_tristate_controller_uas_writedata     (mm_interconnect_0_generic_tristate_controller_uas_writedata),     //                                .writedata
		.generic_tristate_controller_uas_burstcount    (mm_interconnect_0_generic_tristate_controller_uas_burstcount),    //                                .burstcount
		.generic_tristate_controller_uas_byteenable    (mm_interconnect_0_generic_tristate_controller_uas_byteenable),    //                                .byteenable
		.generic_tristate_controller_uas_readdatavalid (mm_interconnect_0_generic_tristate_controller_uas_readdatavalid), //                                .readdatavalid
		.generic_tristate_controller_uas_waitrequest   (mm_interconnect_0_generic_tristate_controller_uas_waitrequest),   //                                .waitrequest
		.generic_tristate_controller_uas_lock          (mm_interconnect_0_generic_tristate_controller_uas_lock),          //                                .lock
		.generic_tristate_controller_uas_debugaccess   (mm_interconnect_0_generic_tristate_controller_uas_debugaccess),   //                                .debugaccess
		.jtag_uart_avalon_jtag_slave_address           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),           //     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),             //                                .write
		.jtag_uart_avalon_jtag_slave_read              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),              //                                .read
		.jtag_uart_avalon_jtag_slave_readdata          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),          //                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),         //                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),       //                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),        //                                .chipselect
		.keyirq_s1_address                             (mm_interconnect_0_keyirq_s1_address),                             //                       keyirq_s1.address
		.keyirq_s1_write                               (mm_interconnect_0_keyirq_s1_write),                               //                                .write
		.keyirq_s1_readdata                            (mm_interconnect_0_keyirq_s1_readdata),                            //                                .readdata
		.keyirq_s1_writedata                           (mm_interconnect_0_keyirq_s1_writedata),                           //                                .writedata
		.keyirq_s1_chipselect                          (mm_interconnect_0_keyirq_s1_chipselect),                          //                                .chipselect
		.keyvalue_s1_address                           (mm_interconnect_0_keyvalue_s1_address),                           //                     keyvalue_s1.address
		.keyvalue_s1_readdata                          (mm_interconnect_0_keyvalue_s1_readdata),                          //                                .readdata
		.lcd_avalon_slave_address                      (mm_interconnect_0_lcd_avalon_slave_address),                      //                lcd_avalon_slave.address
		.lcd_avalon_slave_write                        (mm_interconnect_0_lcd_avalon_slave_write),                        //                                .write
		.lcd_avalon_slave_read                         (mm_interconnect_0_lcd_avalon_slave_read),                         //                                .read
		.lcd_avalon_slave_readdata                     (mm_interconnect_0_lcd_avalon_slave_readdata),                     //                                .readdata
		.lcd_avalon_slave_writedata                    (mm_interconnect_0_lcd_avalon_slave_writedata),                    //                                .writedata
		.lcd_avalon_slave_chipselect                   (mm_interconnect_0_lcd_avalon_slave_chipselect),                   //                                .chipselect
		.sdram_s1_address                              (mm_interconnect_0_sdram_s1_address),                              //                        sdram_s1.address
		.sdram_s1_write                                (mm_interconnect_0_sdram_s1_write),                                //                                .write
		.sdram_s1_read                                 (mm_interconnect_0_sdram_s1_read),                                 //                                .read
		.sdram_s1_readdata                             (mm_interconnect_0_sdram_s1_readdata),                             //                                .readdata
		.sdram_s1_writedata                            (mm_interconnect_0_sdram_s1_writedata),                            //                                .writedata
		.sdram_s1_byteenable                           (mm_interconnect_0_sdram_s1_byteenable),                           //                                .byteenable
		.sdram_s1_readdatavalid                        (mm_interconnect_0_sdram_s1_readdatavalid),                        //                                .readdatavalid
		.sdram_s1_waitrequest                          (mm_interconnect_0_sdram_s1_waitrequest),                          //                                .waitrequest
		.sdram_s1_chipselect                           (mm_interconnect_0_sdram_s1_chipselect),                           //                                .chipselect
		.sysid_control_slave_address                   (mm_interconnect_0_sysid_control_slave_address),                   //             sysid_control_slave.address
		.sysid_control_slave_readdata                  (mm_interconnect_0_sysid_control_slave_readdata),                  //                                .readdata
		.TAS_scl_s1_address                            (mm_interconnect_0_tas_scl_s1_address),                            //                      TAS_scl_s1.address
		.TAS_scl_s1_write                              (mm_interconnect_0_tas_scl_s1_write),                              //                                .write
		.TAS_scl_s1_readdata                           (mm_interconnect_0_tas_scl_s1_readdata),                           //                                .readdata
		.TAS_scl_s1_writedata                          (mm_interconnect_0_tas_scl_s1_writedata),                          //                                .writedata
		.TAS_scl_s1_chipselect                         (mm_interconnect_0_tas_scl_s1_chipselect),                         //                                .chipselect
		.TAS_sda_s1_address                            (mm_interconnect_0_tas_sda_s1_address),                            //                      TAS_sda_s1.address
		.TAS_sda_s1_write                              (mm_interconnect_0_tas_sda_s1_write),                              //                                .write
		.TAS_sda_s1_readdata                           (mm_interconnect_0_tas_sda_s1_readdata),                           //                                .readdata
		.TAS_sda_s1_writedata                          (mm_interconnect_0_tas_sda_s1_writedata),                          //                                .writedata
		.TAS_sda_s1_chipselect                         (mm_interconnect_0_tas_sda_s1_chipselect),                         //                                .chipselect
		.timer0_s1_address                             (mm_interconnect_0_timer0_s1_address),                             //                       timer0_s1.address
		.timer0_s1_write                               (mm_interconnect_0_timer0_s1_write),                               //                                .write
		.timer0_s1_readdata                            (mm_interconnect_0_timer0_s1_readdata),                            //                                .readdata
		.timer0_s1_writedata                           (mm_interconnect_0_timer0_s1_writedata),                           //                                .writedata
		.timer0_s1_chipselect                          (mm_interconnect_0_timer0_s1_chipselect),                          //                                .chipselect
		.touch_irq_s1_address                          (mm_interconnect_0_touch_irq_s1_address),                          //                    touch_irq_s1.address
		.touch_irq_s1_write                            (mm_interconnect_0_touch_irq_s1_write),                            //                                .write
		.touch_irq_s1_readdata                         (mm_interconnect_0_touch_irq_s1_readdata),                         //                                .readdata
		.touch_irq_s1_writedata                        (mm_interconnect_0_touch_irq_s1_writedata),                        //                                .writedata
		.touch_irq_s1_chipselect                       (mm_interconnect_0_touch_irq_s1_chipselect),                       //                                .chipselect
		.toucH_scl_s1_address                          (mm_interconnect_0_touch_scl_s1_address),                          //                    toucH_scl_s1.address
		.toucH_scl_s1_write                            (mm_interconnect_0_touch_scl_s1_write),                            //                                .write
		.toucH_scl_s1_readdata                         (mm_interconnect_0_touch_scl_s1_readdata),                         //                                .readdata
		.toucH_scl_s1_writedata                        (mm_interconnect_0_touch_scl_s1_writedata),                        //                                .writedata
		.toucH_scl_s1_chipselect                       (mm_interconnect_0_touch_scl_s1_chipselect),                       //                                .chipselect
		.touch_sda_s1_address                          (mm_interconnect_0_touch_sda_s1_address),                          //                    touch_sda_s1.address
		.touch_sda_s1_write                            (mm_interconnect_0_touch_sda_s1_write),                            //                                .write
		.touch_sda_s1_readdata                         (mm_interconnect_0_touch_sda_s1_readdata),                         //                                .readdata
		.touch_sda_s1_writedata                        (mm_interconnect_0_touch_sda_s1_writedata),                        //                                .writedata
		.touch_sda_s1_chipselect                       (mm_interconnect_0_touch_sda_s1_chipselect)                        //                                .chipselect
	);

	nios2_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
